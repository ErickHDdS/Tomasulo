library verilog;
use verilog.vl_types.all;
entity pratica3 is
    port(
        clock           : in     vl_logic
    );
end pratica3;
