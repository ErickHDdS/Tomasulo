module IQ(Clock, enableOut, instructionOut, done, disponivel);
  
  input Clock, done, disponivel;
  reg [15:0]PC1[50:0];
  
  reg[15:0] i;

  output reg enableOut;
  output reg[15:0]instructionOut;
  
  initial
	begin 
		i = 0;
		//Fila de Instrucoes:
		//[000]offset [000]Rz [000]Rx [000]Ry [0000] opcode
		PC1[0]=16'b0000110010100000; //ADD R3, R1, R2
      PC1[1]=16'b0001010110010001; //SUB R5, R3, R1
      PC1[2]=16'b0001011001100000; //ADD R5, R4, R6 
      PC1[3]=16'b0001101011000100; //MUL R6, R5,R4 
      PC1[4]=16'b0000101010110100; //MUL R2, R5, R3 
      PC1[5]=16'b0001101011000001; //SUB R6, R5, R4 
      PC1[6]=16'b0001101011010000; //ADD R6, R5, R5 
	end

	always @ (posedge Clock)
	begin
	  	if(disponivel == 1'b1)
		begin
			instructionOut = PC1[i];
			enableOut = 1;
			i = i + 1;
	  end
	end
endmodule