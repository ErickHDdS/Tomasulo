module pratica3(clock);
 input clock;
 
 CDB cdb (clock);
 endmodule