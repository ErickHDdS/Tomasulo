library verilog;
use verilog.vl_types.all;
entity CDB is
    port(
        clock           : in     vl_logic
    );
end CDB;
